`timescale 1ns / 1ps


module vehicle_state(clk, rst_n, state_in, data_in, 